module float_converter(
    input  [31:0] i_int,
    output [30:0] o_float
);

assign o_float = (i_int[31]) ? 31'd0                          : // relu
                 (i_int[30]) ? {(8'd157), i_int[30:8]       } :
                 (i_int[29]) ? {(8'd156), i_int[29:7]       } :
                 (i_int[28]) ? {(8'd155), i_int[28:6]       } :
                 (i_int[27]) ? {(8'd154), i_int[27:5]       } :
                 (i_int[26]) ? {(8'd153), i_int[26:4]       } :
                 (i_int[25]) ? {(8'd152), i_int[25:3]       } :
                 (i_int[24]) ? {(8'd151), i_int[24:2]       } :
                 (i_int[23]) ? {(8'd150), i_int[23:1]       } :
                 (i_int[22]) ? {(8'd149), i_int[22:0]       } :
                 (i_int[21]) ? {(8'd148), i_int[21:0],  1'd0} :
                 (i_int[20]) ? {(8'd147), i_int[20:0],  2'd0} :
                 (i_int[19]) ? {(8'd146), i_int[19:0],  3'd0} :
                 (i_int[18]) ? {(8'd145), i_int[18:0],  4'd0} :
                 (i_int[17]) ? {(8'd144), i_int[17:0],  5'd0} :
                 (i_int[16]) ? {(8'd143), i_int[16:0],  6'd0} :
                 (i_int[15]) ? {(8'd142), i_int[15:0],  7'd0} :
                 (i_int[14]) ? {(8'd141), i_int[14:0],  8'd0} :
                 (i_int[13]) ? {(8'd140), i_int[13:0],  9'd0} :
                 (i_int[12]) ? {(8'd139), i_int[12:0], 10'd0} :
                 (i_int[11]) ? {(8'd138), i_int[11:0], 11'd0} :
                 (i_int[10]) ? {(8'd137), i_int[10:0], 12'd0} :
                 (i_int[9])  ? {(8'd136), i_int[9:0],  13'd0} :
                 (i_int[8])  ? {(8'd135), i_int[8:0],  14'd0} :
                 (i_int[7])  ? {(8'd134), i_int[7:0],  15'd0} :
                 (i_int[6])  ? {(8'd133), i_int[6:0],  16'd0} :
                 (i_int[5])  ? {(8'd132), i_int[5:0],  17'd0} :
                 (i_int[4])  ? {(8'd131), i_int[4:0],  18'd0} :
                 (i_int[3])  ? {(8'd130), i_int[3:0],  19'd0} :
                 (i_int[2])  ? {(8'd129), i_int[2:0],  20'd0} :
                 (i_int[1])  ? {(8'd128), i_int[1:0],  21'd0} :
                 (i_int[0])  ? {(8'd127), i_int[0:0],  22'd0} :
                                                       31'd0;  //zero
endmodule